LPF
V1 N001 0 SINE(0 1e-6 1e4) AC 1
C1 N003 0 2e-11
R1 N002 N001 1e3
R2 N003 N002 500

.control
    define binary(run,index) floor(run/(2^index))-2*floor(run/(2^index+1))
    define wc(nom,tol,index,run,numruns) (run >= numruns) ? nom : (binary(run,index) ? nom*(1+tol) : nom*(1-tol))

    options noacct
    let numruns = 4
  	let run = 0
    let tol = 0.1
    set curplot=new          $ create a new plot
	set scratch=$curplot     $ store its name to 'scratch'
    set color0=white
    let rout1 = unitvec(numruns+1)
    let rout2 = unitvec(numruns+1)
    let cutoff=unitvec(numruns+1)

    dowhile run <= numruns
        alter R1 = wc(1000,0.1,0,run,numruns)
        alter R2 = wc(500,0.1,1,run,numruns)
        show R1 : resistance
        show R2 : resistance

        ac dec 40 1e2 100e6

        meas ac ymax MAX v(N003)
        let v3db = ymax/sqrt(2)
        meas ac cut when v(N003)=v3db fall=last
        let {$scratch}.cutoff[run] = cut

        set run = $&run
		set dt = $curplot
		setplot $scratch

        let vout{$run} = {$dt}.v(N003)
        let rout1[$run] = @r1[resistance]
        let rout2[$run] = @r2[resistance]
        setplot $dt
		let run = run + 1
    end

    *plot db({$scratch}.allv)
    plot {$scratch}.cutoff vs {$scratch}.cout
    setplot $scratch
    print rout1 rout2 cutoff
    wrdata worst $&cutoff

.endc

.end