Sensitivy
V1 N001 0 1
R1 N002 N001 5
R2 0 N002 10
R3 N003 N001 5
R4 0 N003 10

.control
    *op
    sens v(N002, N003)
    print all

.endc

.end