* Resistive partition with different ratios for AC/DC (Print V(2))

vin 1 0 DC 10 sin(0 1 50)
r1  1 2 5K
r2  2 0 5K ac=15k

.control
	shell rm v2
	set appendwrite
	let mc_runs = 5
  	let run = 0
	set curplot=new          $ create a new plot
	set curplottitle=abc
	set scratch=$curplot     $ store its name to 'scratch'
	setplot $scratch         $ make 'scratch' the active plot
	*let vout=unitvec(mc_runs)
	let rout=unitvec(mc_runs)
	
* unif: uniform distribution, deviation relativ to nominal value
* aunif: uniform distribution, deviation absolut
* gauss: Gaussian distribution, deviation relativ to nominal value
* agauss: Gaussian distribution, deviation absolut
* limit: if unif. distributed value >=0 then add +avar to nom, else -avar

	define unif(nom, rvar) (nom + (nom*rvar) * sunif(0))
	define aunif(nom, avar) (nom + avar * sunif(0))
	define gauss(nom, rvar, sig) (nom + (nom*rvar)/sig * sgauss(0))
	define agauss(nom, avar, sig) (nom + avar/sig * sgauss(0))
	define limit(nom, avar) (nom + ((sgauss(0) >= 0) ? avar : -avar))

	dowhile run < mc_runs 
		alter r1 = unif(5k, 0.1)
		alter r2 = gauss(5k, 0.1, 1)
		OP
		show r1 : resistance , r2 : resistance
		print v(2)
		wrdata v2 @r1[resistance] v(2)

		set run = $&run
		set dt = $curplot
		setplot $scratch
		let vout{$run}={$dt}.v(2)
		let rout[run] = @r1[resistance] + @r2[resistance]
		setplot $dt
		let run = run + 1
	end	

	plot {$scratch}.allv
.endc

.END
