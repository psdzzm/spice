* Resistive partition with different ratios for AC/DC (Print V(2))

vin 1 0 DC 10 sin(0 1 50)
r1  1 2 5K
r2  2 0 5K ac=15k

.control
set filetype=ascii
options acct
shell rm v2

let start_r = 5k
let stop_r = 10k
let delta_r = 500
let r_act = start_r
set appendwrite

while r_act le stop_r
	alter r1 r_act
	*TRAN 1m 0.1
	OP
	wrdata v2 v(2)
	let r_act = r_act + delta_r
end

.endc

.END
