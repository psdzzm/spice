LPF
V1 N001 0 SINE(0 1 1e4) AC 1
C1 N002 0 2e-11
R1 N002 N001 1e3

.control
    options noacct
    save all
    let mc_runs = 50
  	let run = 0
    let tol = 0.6
    set curplot=new          $ create a new plot
	set scratch=$curplot     $ store its name to 'scratch'
    set color0=white
    let cout = unitvec(mc_runs)
    let cutoff=unitvec(mc_runs)


    let start_r = @c1[capacitance] * (1 - tol / 2)
    let stop_r = @c1[capacitance] * (1 + tol / 2)

    define stepparam(start_r, stop_r, section, num) (start_r + (stop_r - start_r)/(section - 1) * num)

    dowhile run < mc_runs
        alter C1 = stepparam(start_r, stop_r, mc_runs, run)
        show C1 : capacitance
        ac dec 40 1e2 100e6

        let vdb = db(v(N002))
        meas ac cut when vdb=-3
        let {$scratch}.cutoff[run] = cut

        set run = $&run
		set dt = $curplot
		setplot $scratch

        let vout{$run} = {$dt}.v(N002)
        let cout[$run] = @c1[capacitance]
        setplot $dt
		let run = run + 1
    end

    *plot db({$scratch}.allv)
    plot {$scratch}.cutoff vs {$scratch}.cout
    setplot $scratch
    print cout cutoff
    wrdata step cutoff

.endc

.end