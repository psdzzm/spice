* 2ND-ORDER BUTTERWORTH
*
VS	1	0	AC	1
*
R1	1	2	11.2K
R2	2	3	11.2K
C1	2	out	2000PF
C2	3	0	1000PF
*
* UNITY GAIN AMPLIFIER, RA=OPEN, RB=SHORT
RA	4	0	100MEG
RB	4	xop.3	1
XOP	3 4	out	OPAMP1
*
* SINGLE RC FILTER FOR COMPARISON
R10	1	10	15.9K
C10	10	0	1000PF
*
* OPAMP MACRO MODEL, SINGLE-POLE
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   output
*                   |   |   |
.SUBCKT OPAMP1	     1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* DC GAIN (100K) AND POLE 1 (100HZ)
* GBWP = 10MHz
EGAIN   3 0     1 2     100K
RP1     3       4       1K
CP1     4       0       1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER out 0     4 0     1
ROUT    out       6       10
.ENDS
*
* ANALYSIS
* VIEW RESULTS

.control
	save out 1 10 2 3 4
	options wr_singlescale
	ac dec 40 1 1G
	wrdata ac vdb(out) vdb(1) vdb(10) vdb(2) vdb(3) vdb(4) 
.endc
.end
