LPF
V1 N001 0 DC 1 SINE(0 1 1e4) AC 1
C1 out 0 2e-11
R1 out N001 1e3


.end
