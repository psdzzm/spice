OPAMP3_CMR.CIR - OPAMP MODEL W/ CMR
*
* POWER SUPPLIES
VCC	10	0	DC	+15V
VEE	11	0	DC	-15V
*
* SIGNAL SOURCE
VS	1	0	AC 1
*
XOP	1 1 3  10 11	OPAMP3
RL	3	0	10MEG
*
*
* OPAMP MACRO MODEL (INTERMEDIATE LEVEL WITH CMR)
*
*                IN+ IN- OUT  VCC  VEE
.SUBCKT OPAMP3   1   2   81   101   102
* CMR INPUT
RCM1	1	105	1000MEG
RCM2	2	105	1000MEG
EOS	1 9	POLY(1) 30 100	  0 1
*
Q1	5 9	7	NPN
Q2	6 2	8	NPN
RC1	101	5	95.49
RC2	101	6	95.49
RE1	7	4	43.79
RE2	8	4	43.79
I1	4	102	0.001
*
* OPEN-LOOP GAIN, FIRST POLE AND SLEW RATE
G1	100 10	6 5 0.0104719
RP1	10	100	9.549MEG
CP1	10	100	0.0016667UF
*
* OUTPUT STAGE
EOUT	80 100	10 100	1
RO	80	81	100
*
* CMR DC AND 1ST POLE
GCM	100 30	105 100 1E-11
RCM	30	31	1MEG
LCM	31	100	159
*
* INTERNAL REFERENCE
RREF1	101	103	100K
RREF2	103	102	100K
EREF	100 0	103 0 1
R100	100	0	1MEG
*
.model NPN  NPN(BF=50000)
*
.ENDS
*
* ANALYSIS
.AC 	DEC 	5 1 100MEG
*
* VIEW RESULTS
.PRINT	AC 	V(1)
.PROBE
.END
