TIA
I1 0 N002 SINE(0 1e-6 3e6) AC 1
C1 N002 0 2p
XU1 0 N002 V+ V- out LM6171A/NS
V1 V+ 0 15
V2 V- 0 -15
R1 N002 out 39K

.include LM6171A.txt

.control
    options noacct
    save n001 n002
    let mc_runs = 2
  	let run = 0
    set curplot=new          $ create a new plot
	set scratch=$curplot     $ store its name to 'scratch'
    set color0=white
    let cout = unitvec(mc_runs)
    let cutoff=unitvec(mc_runs)
    setseed 10

    dowhile run < mc_runs
        alter C1 = gauss(2p, 0.1, 1)
        ac dec 40 1e3 100e6

        * plot db(v(N001))
        * plot db(mag(v(N001)))
        meas ac ymax MAX v(N001)
        let v3db = ymax/sqrt(2)
        meas ac cut when v(N001)=v3db fall=last

        let {$scratch}.cutoff[run] = cut

        set run = $&run
		set dt = $curplot
		setplot $scratch

        let vout{$run} = {$dt}.v(N001)
        let cout[$run] = @c1[capacitance]
        setplot $dt
		let run = run + 1
    end

    *plot db({$scratch}.allv)
    setplot $scratch
    print cout cutoff
    wrdata tia cutoff
.endc

C2 out N002 0.7p
.ac oct 40 1e2 100e6

.end
