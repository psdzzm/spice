LPF
V1 N001 0 DC 1 SINE(0 1 1e4) AC 1
C1 out 0 2e-11
R1 out N001 1e3

.control
    SAVE out
    options appendwrite wr_singlescale
    show r : resistance , c : capacitance > list
    OP
    shell rm out
    wrdata out out
    ac dec 40 10 1G
    meas ac ymax MAX v(out)
    meas ac fmax MAX_AT v(out)
    let v3db = ymax/sqrt(2)
    meas ac cut when v(out)=v3db fall=last
    plot vdb(out)
    destroy frequency
    wrdata out fmax cut
.endc

.end

