* D:\74133\OneDrive - University of Edinburgh\Career\Internship\Spice\Spice\rc3.asc
V1 N001 0 SINE(0 1 50) AC 1
R1 out N001 1
C1 out 0 1

.control
	option wr_singlescale
 	op
 	wrdata op all
.endc
 
.end
