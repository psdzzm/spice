TIA
I1 0 N002 SINE(0 1e-6 3e6) AC 1
C1 N002 0 2p
XU1 0 N002 V+ V- out LM6171A/NS
V1 V+ 0 15
V2 V- 0 -15
R1 N002 out 39K
C2 out N002 0.7p
.include lib/aLM6171A
.include lib/escape


.end